* efficiency.cir

.MODEL diode D Is=2e-10 Vj=0.632 Tnom=25

Isolar 0 vsolar 9.07
Dp vsolar 0 diode
Rp vsolar 0 100
Rout vload vsolar 10m

Rload vload 0 {Res}

.OP
.STEP PARAM Res 1n 0.2 .1m
.PRINT I(Isolar) I(Rload) V(vload) V(vsolar)
.MEAS max_eff MAX I(Rload)*V(vload)/(V(vsolar)*I(Isolar))
.MEAS opt_r FIND V(vload)/I(Rload) WHEN I(Rload)*V(vload)/(V(vsolar)*I(Isolar))=max_eff
.END
