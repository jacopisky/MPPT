* cell_test.cir

.LIB cell.cir

X1 vcell 0 PVcell duty={cycle}
Vload vcell 0 DC

.DC Vload 0 0.7 0.01
.STEP PARAM cycle LIST 1 0.9 0.8 0.7 0.6 0.5 0.4 0.3 0.2 0.1
.END
