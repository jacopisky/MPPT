* roc.cir

.LIB cell.cir
.MODEL VDMOS VDMOS(Rg=0.9 Vto=2.33 Rd=1.54m Rs=1.04m Rb=2.46m Kp=242.5 Lambda=0.09 Cgdmin=21p Cgdmax=0.37n A=0.6 Cgs=1.11n Cjo=1.4n M=0.75 Is=12.6p VJ=2.5 N=1.12 TT=3n ksubthres=.1 mfg=Infineon Vds=25 Ron=3.6m Qg=8n)
.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB opamp.cir

* defining voltage meter
.SUBCKT VMETER in+ in- vdd gnd out
R1 in- v- 10k
R2 v- out 10k
R3 in+ v+ 10k
R4 v+ gnd 10k
X1 v+ v- vdd gnd out LM124
.ENDS

* defining not logic port
.SUBCKT NOT in out vdd gnd
M1 out in gnd gnd NMOS
M2 out in vdd vdd PMOS
.ENDS

* defining resistive voltage divider
.SUBCKT DIVIDER in gnd out PARAMS: div=2
.param r2 1Meg
R1 in out {r2*(div-1)}
R2 out gnd {r2}
.ENDS

* modified pv module
Xc1 vcell1 0 PVcell duty=1
Xv1 vcell1 0 vdd 0 vc1 VMETER
Me1 vcell12 ec1 vcell1 vcell1 VDMOS
Mb1 vcell12 nec1 0 0 VDMOS
Rpd1 nec1 0 1k

Xc2 vcell2 vcell12 PVcell duty=0.2
Xv2 vcell2 vcell12 vdd 0 vc2 VMETER
Me2 vcell23 ec2 vcell2 vcell2 VDMOS
Mb2 vcell23 nec2 vcell12 vcell12 VDMOS
Rpd2 nec2 0 1k

Xc3 vcell3 vcell23 PVcell duty=1
Xv3 vcell3 vcell23 vdd 0 vc3 VMETER
Me3 vcell34 ec3 vcell3 vcell3 VDMOS
Mb3 vcell34 nec3 vcell23 vcell23 VDMOS
Rpd3 nec3 0 1k

Xc4 vcell4 vcell34 PVcell duty=1
Xv4 vcell4 vcell34 vdd 0 vc4 VMETER
Me4 vload ec4 vcell4 vcell4 VDMOS
Mb4 vload nec4 vcell34 vcell34 VDMOS
Rpd4 nec4 0 1k

* load
Vload vload 0 DC

* measuring cell's average voltage
* NOTE: ncells needs to be equal to #cells
.param ncells 4
Xsense vload 0 vref DIVIDER div={ncells*1.2}

* comparators
Xref1 vc1 vref vdd 0 ec1 LM124
Xref2 vc2 vref vdd 0 ec2 LM124
Xref3 vc3 vref vdd 0 ec3 LM124
Xref4 vc4 vref vdd 0 ec4 LM124

* NOT logic ports (CMOS)
Xn1 ec1 nec1 vdd 0 NOT
Xn2 ec2 nec2 vdd 0 NOT
Xn3 ec3 nec3 vdd 0 NOT
Xn4 ec4 nec4 vdd 0 NOT

* alimentation of logic network
Vdd vdd 0 10

* analysis requests
.DC Vload 0 2.7 1m
.PRINT V(vc1) V(vc2) V(vc3) V(vc4) V(vref)
.PRINT V(ec1) V(ec2) V(ec3) V(ec4)
.PRINT V(nec1) V(nec2) V(nec3) V(nec4)
.PRINT I(Vload) V(vcell4)
.MEAS Pmax MAX I(Vload)*Vload
.MEAS Impp FIND I(Vload) WHEN I(Vload)*Vload=Pmax
.END
